module fsm(state, odd, even, terminal, pause, restart, clk, rst);

input pause, restart, clk, rst;

output[1:0] state;

output odd, even, terminal;



endmodule